One_inst : One PORT MAP (
		result	 => result_sig
	);
