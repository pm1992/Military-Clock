zbitcont_inst : zbitcont PORT MAP (
		result	 => result_sig
	);
