SixCompare_inst : SixCompare PORT MAP (
		dataa	 => dataa_sig,
		AeB	 => AeB_sig
	);
