ob1_inst : ob1 PORT MAP (
		result	 => result_sig
	);
