Zero4bit_inst : Zero4bit PORT MAP (
		result	 => result_sig
	);
