twocmp_inst : twocmp PORT MAP (
		dataa	 => dataa_sig,
		AeB	 => AeB_sig
	);
