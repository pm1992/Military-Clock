Fast200x_inst : Fast200x PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
