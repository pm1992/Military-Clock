TenKCompare_inst : TenKCompare PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		AeB	 => AeB_sig
	);
