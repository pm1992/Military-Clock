IncSW_inst : IncSW PORT MAP (
		data	 => data_sig,
		eq5	 => eq5_sig
	);
