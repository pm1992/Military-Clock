minmax_inst : minmax PORT MAP (
		dataa	 => dataa_sig,
		AlB	 => AlB_sig
	);
