Fourbit1_inst : Fourbit1 PORT MAP (
		result	 => result_sig
	);
