Zero_inst : Zero PORT MAP (
		result	 => result_sig
	);
