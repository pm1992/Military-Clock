FourCounter_inst : FourCounter PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
