FiveKCounter_inst : FiveKCounter PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
